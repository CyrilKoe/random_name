package types_pkg;
    
    typedef enum bit { EVEN=0, ODD=1 } e_parity_mode;
    typedef enum bit { LSB, MSB } e_parity_bit_choice;
    
endpackage: types_pkg
